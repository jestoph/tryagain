---------------------------------------------------------------------------
-- single_cycle_core.vhd - A Single-Cycle Processor Implementation
--
-- Notes : 
--
-- See single_cycle_core.pdf for the block diagram of this single
-- cycle processor core.
--
-- Instruction Set Architecture (ISA) for the single-cycle-core:
--   Each instruction is 16-bit wide, with four 4-bit fields.
--
--     noop      
--        # no operation or to signal end of program
--        # format:  | opcode = 0 |  0   |  0   |   0    | 
--
--     load  rt, rs, offset     
--        # load data at memory location (rs + offset) into rt
--        # format:  | opcode = 1 |  rs  |  rt  | offset |
--
--     store rt, rs, offset
--        # store data rt into memory location (rs + offset)
--        # format:  | opcode = 3 |  rs  |  rt  | offset |
--
--     add   rd, rs, rt
--        # rd <- rs + rt
--        # format:  | opcode = 8 |  rs  |  rt  |   rd   |
--
--
-- Copyright (C) 2006 by Lih Wen Koh (lwkoh@cse.unsw.edu.au)
-- All Rights Reserved. 
--
-- The single-cycle processor core is provided AS IS, with no warranty of 
-- any kind, express or implied. The user of the program accepts full 
-- responsibility for the application of the program and the use of any 
-- results. This work may be downloaded, compiled, executed, copied, and 
-- modified solely for nonprofit, educational, noncommercial research, and 
-- noncommercial scholarship purposes provided that this notice in its 
-- entirety accompanies all copies. Copies of the modified software can be 
-- delivered to persons who use it solely for nonprofit, educational, 
-- noncommercial research, and noncommercial scholarship purposes provided 
-- that this notice in its entirety accompanies all copies.
--
---------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity single_cycle_core is
    port ( reset  : in  std_logic;
           clk    : in  std_logic;
           clk_pc  : in std_logic           );
end single_cycle_core;

architecture structural of single_cycle_core is

component program_counter is
    port ( reset    : in  std_logic;
           clk      : in  std_logic;
           addr_in  : in  std_logic_vector(11 downto 0);
           addr_out : out std_logic_vector(11 downto 0) );
end component;

component instruction_memory is
    port ( reset    : in  std_logic;
           clk      : in  std_logic;
           addr_in  : in  std_logic_vector(11 downto 0);
           insn_out : out std_logic_vector(15 downto 0) );
end component;

component sign_extend_4to16 is
    port ( data_in  : in  std_logic_vector(3 downto 0);
           data_out : out std_logic_vector(15 downto 0) );
end component;

component sign_extend_4to12 is
    port ( data_in  : in  std_logic_vector(3 downto 0);
           data_out : out std_logic_vector(11 downto 0) );
end component;

component mux_2to1_4b is
    port ( mux_select : in  std_logic;
           data_a     : in  std_logic_vector(3 downto 0);
           data_b     : in  std_logic_vector(3 downto 0);
           data_out   : out std_logic_vector(3 downto 0) );
end component;

component mux_2to1_12b is
    port ( mux_select : in  std_logic;
           data_a     : in  std_logic_vector(11 downto 0);
           data_b     : in  std_logic_vector(11 downto 0);
           data_out   : out std_logic_vector(11 downto 0) );
end component;

component mux_2to1_16b is
    port ( mux_select : in  std_logic;
           data_a     : in  std_logic_vector(15 downto 0);
           data_b     : in  std_logic_vector(15 downto 0);
           data_out   : out std_logic_vector(15 downto 0) );
end component;

component control_unit is
    port ( opcode     : in  std_logic_vector(3 downto 0);
           reg_dst    : out std_logic;
           reg_write  : out std_logic;
           alu_src    : out std_logic;
           alu_op	  : out std_logic_vector(2 downto 0);
           mem_write  : out std_logic;
           do_jmp     : out std_logic;
           do_not_jmp : out std_logic;
           do_slt     : out std_logic;
           byte_addr  : out std_logic;
           b_type     : out std_logic;
           b_insn     : out std_logic;
           mem_read   : out std_logic;
           do_branch  : in  std_logic;
           do_pc_offset : out std_logic;
           mem_to_reg : out std_logic );
end component;

component register_file is
    port ( reset           : in  std_logic;
           clk             : in  std_logic;
           read_register_a : in  std_logic_vector(3 downto 0);
           read_register_b : in  std_logic_vector(3 downto 0);
           write_enable    : in  std_logic;
           write_register  : in  std_logic_vector(3 downto 0);
           write_data      : in  std_logic_vector(15 downto 0);
           read_data_a     : out std_logic_vector(15 downto 0);
           read_data_b     : out std_logic_vector(15 downto 0) );
end component;

component adder_4b is
    port ( src_a     : in  std_logic_vector(3 downto 0);
           src_b     : in  std_logic_vector(3 downto 0);
           sum       : out std_logic_vector(3 downto 0);
           carry_out : out std_logic );
end component;

component alu_16b is
    port ( src_a     : in  std_logic_vector(15 downto 0);
           src_b     : in  std_logic_vector(15 downto 0);
           alu_out   : out std_logic_vector(15 downto 0);
           alu_op	 : in  std_logic_vector(2 downto 0);
           do_slt    : in  std_logic;
           carry_out : out std_logic );
end component;

component data_memory is
    port ( reset        : in  std_logic;
           clk          : in  std_logic;
           write_enable : in  std_logic;
           read_enable  : in  std_logic;
           write_data   : in  std_logic_vector(15 downto 0);
           byte_addr	   : in  std_logic;
           addr_in      : in  std_logic_vector(11 downto 0);
           data_out     : out std_logic_vector(15 downto 0) );
end component;

component branch_cmp is
    port ( b_type       : in  std_logic; -- 1 for beq
           b_insn       : in  std_logic; -- 1 for b instruction
           src_a        : in  std_logic_vector(15 downto 0);
           src_b        : in  std_logic_vector(15 downto 0);
           do_branch    : out std_logic); -- 1 if doing branch
end component;

component adder_12b is
    port ( src_a     : in  std_logic_vector(11 downto 0);
           src_b     : in  std_logic_vector(11 downto 0);
           sum       : out std_logic_vector(11 downto 0);
           carry_in  : in  std_logic;
           carry_out : out std_logic );
end component;

--------------------------------------------------------------
-- pipeline registers
--
--------------------------------------------------------------

component generic_register is
    port ( reset        : in  std_logic;
           clk          : in  std_logic;
           data_out		: out std_logic_vector(15 downto 0);
           data_in     	: in  std_logic_vector(15 downto 0));
end component;


signal sig_next_pc              : std_logic_vector(11 downto 0);
signal sig_curr_pc              : std_logic_vector(11 downto 0);
signal sig_one_4b               : std_logic_vector(3 downto 0);
signal sig_one_12b              : std_logic_vector(11 downto 0);
signal sig_pc_carry_out         : std_logic;
signal sig_insn                 : std_logic_vector(15 downto 0);
signal sig_sign_extended_offset : std_logic_vector(15 downto 0);
signal sig_reg_dst              : std_logic;
signal sig_reg_write            : std_logic;
signal sig_alu_src              : std_logic;
signal sig_mem_write            : std_logic;
signal sig_mem_to_reg           : std_logic;
signal sig_write_register       : std_logic_vector(3 downto 0);
signal sig_write_data           : std_logic_vector(15 downto 0);
signal sig_read_data_a          : std_logic_vector(15 downto 0);
signal sig_read_data_b          : std_logic_vector(15 downto 0);
signal sig_alu_src_b            : std_logic_vector(15 downto 0);
signal sig_alu_result           : std_logic_vector(15 downto 0); 
signal sig_alu_carry_out        : std_logic;
signal sig_data_mem_out         : std_logic_vector(15 downto 0);
signal sig_alu_op			        : std_logic_vector(2 downto 0);
signal sig_do_slt               : std_logic;
signal sig_byte_addr            : std_logic;
signal sig_mem_read             : std_logic;
signal sig_b_type               : std_logic;
signal sig_b_insn               : std_logic;

-- The following are added to allow for modifications to the pc
-- ie for branching and jumping.
-- When jumping (signaled by sig_do_jmp=1) we read the address from
-- the immediate that is within the instruction itself
-- When branching we still read the address from the instruction 
-- immediate, but in this case it is a 4-bit value so must be sign extended 
-- NOTE! The instruction memory is limited to 2^12 addresses for 
-- convenience.


signal sig_do_branch            : std_logic;
signal sig_do_jmp               : std_logic;
signal sig_curr_pc_or_branch    : std_logic_vector(11 downto 0);
signal sig_branch_offset        : std_logic_vector(11 downto 0);
signal sig_z_12b                : std_logic_vector(11 downto 0);
signal sig_jump_or_branch_addr  : std_logic_vector(11 downto 0);
signal sig_do_pc_offset         : std_logic;
signal sig_pc_or_jmp            : std_logic_vector(11 downto 0);
signal sig_z_or_branch          : std_logic_vector(11 downto 0);
signal sig_one_or_branch        : std_logic_vector(11 downto 0);
signal sig_do_not_jmp           : std_logic;

-------------------------------------------
-- Pipeline signals
-- 
-------------------------------------------
signal sig_next_pc_if           : std_logic_vector(11 downto 0);
signal sig_next_pc_id           : std_logic_vector(11 downto 0);
signal sig_insn_if              : std_logic_vector(15 downto 0);

begin

    sig_one_4b <= "0001";
	 sig_one_12b <= "000000000001";
    sig_z_12b <= "000000000000";
    

    pc : program_counter
    port map ( reset    => reset,
               clk      => clk,
               addr_in  => sig_next_pc,
               addr_out => sig_curr_pc ); 

    -- We need to sign extend because a branch encodes the address in an immediate
    branch_extend : sign_extend_4to12 
    port map ( data_in  => sig_insn(3 downto 0),
               data_out => sig_branch_offset );

    -- Choose whether we're branching or not
    -- or from an immediate (j)
    pc_mux_bjmp : mux_2to1_12b 
    port map ( mux_select => sig_do_branch,
               data_a     => sig_z_12b, -- or we don't branch
               data_b     => sig_branch_offset, -- Branch has address encoded in last nibble
               data_out   => sig_one_or_branch);
    

    -- Choose whether we go to an absolute jump or not 
    pc_mux_offset : mux_2to1_12b 
    port map ( mux_select => sig_do_jmp,
               data_a     => sig_curr_pc, --or not jump
               data_b     => sig_insn(11 downto 0), --we can jump
               data_out   => sig_pc_or_jmp);

    next_pc : adder_12b 
    port map ( src_a     => sig_pc_or_jmp, 
               src_b     => sig_one_or_branch,
               sum       => sig_next_pc,   
               carry_in  => sig_do_not_jmp,
               carry_out => sig_pc_carry_out );
    
    insn_mem : instruction_memory 
    port map ( reset    => reset,
               clk      => clk,
               addr_in  => sig_next_pc,
               insn_out => sig_insn_if );

    sign_extend : sign_extend_4to16 
    port map ( data_in  => sig_insn(3 downto 0),
               data_out => sig_sign_extended_offset );

    ctrl_unit : control_unit 
    port map ( opcode     => sig_insn(15 downto 12),
               reg_dst    => sig_reg_dst,
               reg_write  => sig_reg_write,
               alu_src    => sig_alu_src,
               mem_write  => sig_mem_write,
               mem_read   => sig_mem_read,
               mem_to_reg => sig_mem_to_reg,
               do_jmp     => sig_do_jmp,
               do_not_jmp => sig_do_not_jmp,
               do_slt     => sig_do_slt,
               byte_addr  => sig_byte_addr,
               b_type     => sig_b_type,
               b_insn     => sig_b_insn,
               do_branch  => sig_do_branch,
               do_pc_offset => sig_do_pc_offset,
			   alu_op	  => sig_alu_op);

    mux_reg_dst : mux_2to1_4b 
    port map ( mux_select => sig_reg_dst,
               data_a     => sig_insn(7 downto 4),
               data_b     => sig_insn(3 downto 0),
               data_out   => sig_write_register );

    reg_file : register_file 
    port map ( reset           => reset, 
               clk             => clk,
               read_register_a => sig_insn(11 downto 8),
               read_register_b => sig_insn(7 downto 4),
               write_enable    => sig_reg_write,
               write_register  => sig_write_register,
               write_data      => sig_write_data,
               read_data_a     => sig_read_data_a,
               read_data_b     => sig_read_data_b );
               
    reg_cmp   : branch_cmp
    port map ( b_type     => sig_b_type,
               b_insn     => sig_b_insn,
               src_a      => sig_read_data_a,
               src_b      => sig_read_data_b,
               do_branch  => sig_do_branch);
    
    mux_alu_src : mux_2to1_16b 
    port map ( mux_select => sig_alu_src,
               data_a     => sig_read_data_b,
               data_b     => sig_sign_extended_offset,
               data_out   => sig_alu_src_b );

    alu : alu_16b 
    port map ( src_a      => sig_read_data_a,
               src_b      => sig_alu_src_b,
               alu_out    => sig_alu_result,
			   alu_op 	  => sig_alu_op,
               do_slt     => sig_do_slt,
               carry_out  => sig_alu_carry_out );

    data_mem : data_memory 
    port map ( reset        => reset,
               clk          => clk,
               write_enable => sig_mem_write,
               read_enable  => sig_mem_read,
               write_data   => sig_read_data_b,
               byte_addr	=> sig_byte_addr,
               addr_in      => sig_alu_result(11 downto 0),
               data_out     => sig_data_mem_out );
               
    mux_mem_to_reg : mux_2to1_16b 
    port map ( mux_select => sig_mem_to_reg,
               data_a     => sig_alu_result,
               data_b     => sig_data_mem_out,
               data_out   => sig_write_data );

----------------------------------------------------
-- Pipeline registers
--
----------------------------------------------------

   register_if_id   : generic_register
    port map(  reset       => reset,
               clk         => clk,
               data_out	   => sig_insn,
               data_in     => sig_insn_if);

end structural;
